/*Approx int16*/
module mul_unit (out, a, b);
	output [31:0] out;
        input [15:0] a;
        input [15:0] b;

 	wire [15:0] a_magnitude; 
 	wire [15:0] b_magnitude; 
 	wire [31:0] mult_out; 
 	wire [31:0] mult_out_2c; 
 	wire sign_m;
  	wire [15:0] wire_pp1; 
  	wire [15:0] wire_pp2; 
  	wire [15:0] wire_pp3; 
  	wire [15:0] wire_pp4; 

	
        assign a_magnitude = (a[15])? (~a+1) : a;
	assign b_magnitude = (b[15])? (~b+1) : b;
	assign sign_m = a[15]^b[15];
	assign mult_out = { 8'b0, wire_pp2, 8'b0} + {8'b0, wire_pp3, 8'b0} + {wire_pp4, wire_pp1};
	assign mult_out_2c = (sign_m)? ((~mult_out)+1) : mult_out;
	assign out = mult_out_2c;
	
mult8x8 u_mult8_pp1(
.a          ( a_magnitude[7:0] ),
.b          ( b_magnitude[7:0] ),
.out        ( wire_pp1 )
);

mult8x8 u_mult8_pp2(
.a          ( a_magnitude[15:8] ),
.b          ( b_magnitude[7:0] ),
.out        ( wire_pp2 )
);

mult8x8 u_mult8_pp3(
.a          ( a_magnitude[7:0] ),
.b          ( b_magnitude[15:8] ),
.out        ( wire_pp3 )
);

mult8x8 u_mult8_pp4(
.a          ( a_magnitude[15:8] ),
.b          ( b_magnitude[15:8] ),
.out        ( wire_pp4 )
);

endmodule


