module mult8x8_inference (
  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
  y16, y15, y14, y13, y12, y11, y10, y9, y8, y7, y6, y5, y4, y3, y2, y1
);
input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15;
output y16, y15, y14, y13, y12, y11, y10, y9, y8, y7, y6, y5, y4, y3, y2, y1;
wire w161, w162, w163, w164, w165, w166, w167, w168, w169, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w151, w152, w153, w154, w155, w156, w157, w158, w159, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w141, w142, w143, w144, w145, w146, w147, w148, w149, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w131, w132, w133, w134, w135, w136, w137, w138, w139, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w121, w122, w123, w124, w125, w126, w127, w128, w129, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w111, w112, w113, w114, w115, w116, w117, w118, w119, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w101, w102, w103, w104, w105, w106, w107, w108, w109, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w91, w92, w93, w94, w95, w96, w97, w98, w99, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w81, w82, w83, w84, w85, w86, w87, w88, w89, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w71, w72, w73, w74, w75, w76, w77, w78, w79, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w61, w62, w63, w64, w65, w66, w67, w68, w69, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w51, w52, w53, w54, w55, w56, w57, w58, w59, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w41, w42, w43, w44, w45, w46, w47, w48, w49, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w31, w32, w33, w34, w35, w36, w37, w38, w39, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w21, w22, w23, w24, w25, w26, w27, w28, w29, w210, w211, w212, w213, w214, w215, w216, w217, w11, w12, w13, w14, w15;
assign w161 = x0 ? w163 : w162;
assign w162 = 0;
assign w163 = x8 ? w165 : w164;
assign w164 = 0;
assign w165 = x1 ? w167 : w166;
assign w166 = x9 ? w169 : w168;
assign w167 = x9 ? w1611 : w1610;
assign w168 = x2 ? w1613 : w1612;
assign w169 = x2 ? w1615 : w1614;
assign w1610 = x10 ? w1617 : w1616;
assign w1611 = 1;
assign w1612 = 0;
assign w1613 = x10 ? w1619 : w1618;
assign w1614 = x10 ? w1621 : w1620;
assign w1615 = x3 ? w1623 : w1622;
assign w1616 = x2 ? w1625 : w1624;
assign w1617 = x2 ? w1627 : w1626;
assign w1618 = 0;
assign w1619 = x3 ? w1629 : w1628;
assign w1620 = x3 ? w1631 : w1630;
assign w1621 = x3 ? w1633 : w1632;
assign w1622 = x10 ? w1635 : w1634;
assign w1623 = 1;
assign w1624 = x11 ? w1637 : w1636;
assign w1625 = x11 ? w1639 : w1638;
assign w1626 = x3 ? w1641 : w1640;
assign w1627 = 1;
assign w1628 = 0;
assign w1629 = x11 ? w1643 : w1642;
assign w1630 = 0;
assign w1631 = x11 ? w1645 : w1644;
assign w1632 = x11 ? w1647 : w1646;
assign w1633 = 1;
assign w1634 = x11 ? w1649 : w1648;
assign w1635 = 1;
assign w1636 = 0;
assign w1637 = x3 ? w1651 : w1650;
assign w1638 = x3 ? w1653 : w1652;
assign w1639 = 1;
assign w1640 = x11 ? w1655 : w1654;
assign w1641 = 1;
assign w1642 = 0;
assign w1643 = x4 ? w1657 : w1656;
assign w1644 = 0;
assign w1645 = x4 ? w1659 : w1658;
assign w1646 = 0;
assign w1647 = x4 ? w1661 : w1660;
assign w1648 = x4 ? w1663 : w1662;
assign w1649 = 1;
assign w1650 = 0;
assign w1651 = x12 ? w1665 : w1664;
assign w1652 = x12 ? w1667 : w1666;
assign w1653 = x12 ? w1669 : w1668;
assign w1654 = x12 ? w1671 : w1670;
assign w1655 = 1;
assign w1656 = x12 ? w1673 : w1672;
assign w1657 = 1;
assign w1658 = 0;
assign w1659 = 1;
assign w1660 = x5 ? w1675 : w1674;
assign w1661 = 1;
assign w1662 = x12 ? w1677 : w1676;
assign w1663 = 1;
assign w1664 = 0;
assign w1665 = 1;
assign w1666 = 0;
assign w1667 = x4 ? w1679 : w1678;
assign w1668 = 0;
assign w1669 = 1;
assign w1670 = x4 ? w1681 : w1680;
assign w1671 = 1;
assign w1672 = 0;
assign w1673 = 1;
assign w1674 = 0;
assign w1675 = 1;
assign w1676 = 0;
assign w1677 = 1;
assign w1678 = 0;
assign w1679 = 1;
assign w1680 = 0;
assign w1681 = 1;
assign w151 = x0 ? w153 : w152;
assign w152 = x1 ? w155 : w154;
assign w153 = x8 ? w157 : w156;
assign w154 = 0;
assign w155 = x8 ? w159 : w158;
assign w156 = x9 ? w1511 : w1510;
assign w157 = x1 ? w1513 : w1512;
assign w158 = 0;
assign w159 = x2 ? w1515 : w1514;
assign w1510 = 0;
assign w1511 = x10 ? w1517 : w1516;
assign w1512 = x9 ? w1519 : w1518;
assign w1513 = x9 ? w1521 : w1520;
assign w1514 = x9 ? w1523 : w1522;
assign w1515 = x9 ? w1525 : w1524;
assign w1516 = x1 ? w1527 : w1526;
assign w1517 = x1 ? w1529 : w1528;
assign w1518 = 1;
assign w1519 = x2 ? w1531 : w1530;
assign w1520 = x10 ? w1533 : w1532;
assign w1521 = x2 ? w1535 : w1534;
assign w1522 = 0;
assign w1523 = x3 ? w1537 : w1536;
assign w1524 = x10 ? w1539 : w1538;
assign w1525 = 1;
assign w1526 = 0;
assign w1527 = x11 ? w1541 : w1540;
assign w1528 = x2 ? w1543 : w1542;
assign w1529 = 1;
assign w1530 = x10 ? w1545 : w1544;
assign w1531 = 0;
assign w1532 = x2 ? w1547 : w1546;
assign w1533 = 0;
assign w1534 = x10 ? w1549 : w1548;
assign w1535 = x10 ? w1551 : w1550;
assign w1536 = x10 ? w1553 : w1552;
assign w1537 = 1;
assign w1538 = x3 ? w1555 : w1554;
assign w1539 = 1;
assign w1540 = x2 ? w1557 : w1556;
assign w1541 = 1;
assign w1542 = x11 ? w1559 : w1558;
assign w1543 = 1;
assign w1544 = 1;
assign w1545 = x3 ? w1561 : w1560;
assign w1546 = 1;
assign w1547 = x11 ? w1563 : w1562;
assign w1548 = 0;
assign w1549 = x3 ? w1565 : w1564;
assign w1550 = x11 ? w1567 : w1566;
assign w1551 = 1;
assign w1552 = 0;
assign w1553 = 1;
assign w1554 = 0;
assign w1555 = 1;
assign w1556 = 0;
assign w1557 = 1;
assign w1558 = 0;
assign w1559 = 1;
assign w1560 = 1;
assign w1561 = 0;
assign w1562 = 1;
assign w1563 = 0;
assign w1564 = 0;
assign w1565 = 1;
assign w1566 = 0;
assign w1567 = 1;
assign w141 = x0 ? w143 : w142;
assign w142 = x1 ? w145 : w144;
assign w143 = x9 ? w147 : w146;
assign w144 = x2 ? w149 : w148;
assign w145 = x8 ? w1411 : w1410;
assign w146 = x10 ? w1413 : w1412;
assign w147 = x10 ? w1415 : w1414;
assign w148 = 0;
assign w149 = x8 ? w1417 : w1416;
assign w1410 = x9 ? w1419 : w1418;
assign w1411 = x2 ? w1421 : w1420;
assign w1412 = x8 ? w1423 : w1422;
assign w1413 = x11 ? w1425 : w1424;
assign w1414 = x2 ? w1427 : w1426;
assign w1415 = x1 ? w1429 : w1428;
assign w1416 = 0;
assign w1417 = x3 ? w1431 : w1430;
assign w1418 = 0;
assign w1419 = x2 ? w1433 : w1432;
assign w1420 = x9 ? w1435 : w1434;
assign w1421 = x9 ? w1437 : w1436;
assign w1422 = 0;
assign w1423 = x1 ? w1439 : w1438;
assign w1424 = x2 ? w1441 : w1440;
assign w1425 = x2 ? w1443 : w1442;
assign w1426 = x1 ? w1445 : w1444;
assign w1427 = x11 ? w1447 : w1446;
assign w1428 = x11 ? w1449 : w1448;
assign w1429 = x2 ? w1451 : w1450;
assign w1430 = x9 ? w1453 : w1452;
assign w1431 = 1;
assign w1432 = x10 ? w1455 : w1454;
assign w1433 = 1;
assign w1434 = 1;
assign w1435 = x3 ? w1457 : w1456;
assign w1436 = x10 ? w1459 : w1458;
assign w1437 = x3 ? w1461 : w1460;
assign w1438 = x2 ? w1463 : w1462;
assign w1439 = x2 ? w1465 : w1464;
assign w1440 = 0;
assign w1441 = x3 ? w1467 : w1466;
assign w1442 = x8 ? w1469 : w1468;
assign w1443 = 1;
assign w1444 = 1;
assign w1445 = x8 ? w1471 : w1470;
assign w1446 = x3 ? w1473 : w1472;
assign w1447 = x1 ? w1475 : w1474;
assign w1448 = x2 ? w1477 : w1476;
assign w1449 = 0;
assign w1450 = 0;
assign w1451 = x11 ? w1479 : w1478;
assign w1452 = 0;
assign w1453 = 1;
assign w1454 = 0;
assign w1455 = 1;
assign w1456 = 1;
assign w1457 = 0;
assign w1458 = 1;
assign w1459 = 0;
assign w1460 = 0;
assign w1461 = 1;
assign w1462 = 0;
assign w1463 = 1;
assign w1464 = 1;
assign w1465 = 0;
assign w1466 = 0;
assign w1467 = 1;
assign w1468 = 1;
assign w1469 = x1 ? w1481 : w1480;
assign w1470 = x11 ? w1483 : w1482;
assign w1471 = 1;
assign w1472 = 1;
assign w1473 = 0;
assign w1474 = x8 ? w1485 : w1484;
assign w1475 = 0;
assign w1476 = 1;
assign w1477 = 0;
assign w1478 = 0;
assign w1479 = 1;
assign w1480 = 1;
assign w1481 = 0;
assign w1482 = 1;
assign w1483 = 0;
assign w1484 = 1;
assign w1485 = 0;
assign w131 = x0 ? w133 : w132;
assign w132 = x1 ? w135 : w134;
assign w133 = x10 ? w137 : w136;
assign w134 = x2 ? w139 : w138;
assign w135 = x9 ? w1311 : w1310;
assign w136 = x11 ? w1313 : w1312;
assign w137 = x11 ? w1315 : w1314;
assign w138 = x3 ? w1317 : w1316;
assign w139 = x8 ? w1319 : w1318;
assign w1310 = x10 ? w1321 : w1320;
assign w1311 = x3 ? w1323 : w1322;
assign w1312 = x8 ? w1325 : w1324;
assign w1313 = x12 ? w1327 : w1326;
assign w1314 = x3 ? w1329 : w1328;
assign w1315 = x1 ? w1331 : w1330;
assign w1316 = 0;
assign w1317 = x8 ? w1333 : w1332;
assign w1318 = x9 ? w1335 : w1334;
assign w1319 = x3 ? w1337 : w1336;
assign w1320 = x8 ? w1339 : w1338;
assign w1321 = x11 ? w1341 : w1340;
assign w1322 = x10 ? w1343 : w1342;
assign w1323 = x10 ? w1345 : w1344;
assign w1324 = x9 ? w1347 : w1346;
assign w1325 = x2 ? w1349 : w1348;
assign w1326 = x3 ? w1351 : w1350;
assign w1327 = x8 ? w1353 : w1352;
assign w1328 = 1;
assign w1329 = x12 ? w1355 : w1354;
assign w1330 = x3 ? w1357 : w1356;
assign w1331 = x12 ? w1359 : w1358;
assign w1332 = 0;
assign w1333 = x4 ? w1361 : w1360;
assign w1334 = 0;
assign w1335 = x3 ? w1363 : w1362;
assign w1336 = x9 ? w1365 : w1364;
assign w1337 = 0;
assign w1338 = 0;
assign w1339 = x2 ? w1367 : w1366;
assign w1340 = x3 ? w1369 : w1368;
assign w1341 = 1;
assign w1342 = 1;
assign w1343 = x4 ? w1371 : w1370;
assign w1344 = x11 ? w1373 : w1372;
assign w1345 = x11 ? w1375 : w1374;
assign w1346 = 0;
assign w1347 = x1 ? w1377 : w1376;
assign w1348 = x3 ? w1379 : w1378;
assign w1349 = x3 ? w1381 : w1380;
assign w1350 = 0;
assign w1351 = 1;
assign w1352 = 1;
assign w1353 = x3 ? w1383 : w1382;
assign w1354 = x4 ? w1385 : w1384;
assign w1355 = 0;
assign w1356 = x4 ? w1387 : w1386;
assign w1357 = x9 ? w1389 : w1388;
assign w1358 = 0;
assign w1359 = x3 ? w1391 : w1390;
assign w1360 = 0;
assign w1361 = 1;
assign w1362 = 0;
assign w1363 = 1;
assign w1364 = 1;
assign w1365 = 0;
assign w1366 = 0;
assign w1367 = 1;
assign w1368 = 0;
assign w1369 = 1;
assign w1370 = 1;
assign w1371 = 0;
assign w1372 = 1;
assign w1373 = 0;
assign w1374 = 0;
assign w1375 = 1;
assign w1376 = 0;
assign w1377 = 1;
assign w1378 = 0;
assign w1379 = 1;
assign w1380 = 1;
assign w1381 = 0;
assign w1382 = 0;
assign w1383 = 1;
assign w1384 = 1;
assign w1385 = 0;
assign w1386 = 1;
assign w1387 = 0;
assign w1388 = 0;
assign w1389 = 1;
assign w1390 = 0;
assign w1391 = 1;
assign w121 = x0 ? w123 : w122;
assign w122 = x1 ? w125 : w124;
assign w123 = x11 ? w127 : w126;
assign w124 = x2 ? w129 : w128;
assign w125 = x10 ? w1211 : w1210;
assign w126 = x12 ? w1213 : w1212;
assign w127 = x12 ? w1215 : w1214;
assign w128 = x3 ? w1217 : w1216;
assign w129 = x9 ? w1219 : w1218;
assign w1210 = x11 ? w1221 : w1220;
assign w1211 = x11 ? w1223 : w1222;
assign w1212 = x8 ? w1225 : w1224;
assign w1213 = x13 ? w1227 : w1226;
assign w1214 = x4 ? w1229 : w1228;
assign w1215 = 0;
assign w1216 = x4 ? w1231 : w1230;
assign w1217 = x8 ? w1233 : w1232;
assign w1218 = x10 ? w1235 : w1234;
assign w1219 = x4 ? w1237 : w1236;
assign w1220 = x8 ? w1239 : w1238;
assign w1221 = x12 ? w1241 : w1240;
assign w1222 = x4 ? w1243 : w1242;
assign w1223 = x2 ? w1245 : w1244;
assign w1224 = x9 ? w1247 : w1246;
assign w1225 = x3 ? w1249 : w1248;
assign w1226 = x4 ? w1251 : w1250;
assign w1227 = x4 ? w1253 : w1252;
assign w1228 = 1;
assign w1229 = x13 ? w1255 : w1254;
assign w1230 = 0;
assign w1231 = x8 ? w1257 : w1256;
assign w1232 = x9 ? w1259 : w1258;
assign w1233 = x4 ? w1261 : w1260;
assign w1234 = 0;
assign w1235 = x4 ? w1263 : w1262;
assign w1236 = x10 ? w1265 : w1264;
assign w1237 = 0;
assign w1238 = 0;
assign w1239 = x3 ? w1267 : w1266;
assign w1240 = x4 ? w1269 : w1268;
assign w1241 = 1;
assign w1242 = 1;
assign w1243 = x12 ? w1271 : w1270;
assign w1244 = 0;
assign w1245 = x12 ? w1273 : w1272;
assign w1246 = 0;
assign w1247 = x2 ? w1275 : w1274;
assign w1248 = x4 ? w1277 : w1276;
assign w1249 = x4 ? w1279 : w1278;
assign w1250 = 0;
assign w1251 = 1;
assign w1252 = x8 ? w1281 : w1280;
assign w1253 = 1;
assign w1254 = 1;
assign w1255 = 0;
assign w1256 = 0;
assign w1257 = 1;
assign w1258 = 0;
assign w1259 = 1;
assign w1260 = 1;
assign w1261 = 0;
assign w1262 = 0;
assign w1263 = 1;
assign w1264 = 1;
assign w1265 = 0;
assign w1266 = 0;
assign w1267 = 1;
assign w1268 = 0;
assign w1269 = 1;
assign w1270 = 1;
assign w1271 = 0;
assign w1272 = 0;
assign w1273 = 1;
assign w1274 = 0;
assign w1275 = 1;
assign w1276 = 0;
assign w1277 = 1;
assign w1278 = 1;
assign w1279 = 0;
assign w1280 = 1;
assign w1281 = 0;
assign w111 = x0 ? w113 : w112;
assign w112 = x1 ? w115 : w114;
assign w113 = x12 ? w117 : w116;
assign w114 = x2 ? w119 : w118;
assign w115 = x11 ? w1111 : w1110;
assign w116 = x13 ? w1113 : w1112;
assign w117 = x13 ? w1115 : w1114;
assign w118 = x3 ? w1117 : w1116;
assign w119 = x10 ? w1119 : w1118;
assign w1110 = x12 ? w1121 : w1120;
assign w1111 = x12 ? w1123 : w1122;
assign w1112 = x8 ? w1125 : w1124;
assign w1113 = x14 ? w1127 : w1126;
assign w1114 = x5 ? w1129 : w1128;
assign w1115 = x5 ? w1131 : w1130;
assign w1116 = x4 ? w1133 : w1132;
assign w1117 = x9 ? w1135 : w1134;
assign w1118 = x11 ? w1137 : w1136;
assign w1119 = x11 ? w1139 : w1138;
assign w1120 = x8 ? w1141 : w1140;
assign w1121 = x13 ? w1143 : w1142;
assign w1122 = x5 ? w1145 : w1144;
assign w1123 = x5 ? w1147 : w1146;
assign w1124 = x9 ? w1149 : w1148;
assign w1125 = x4 ? w1151 : w1150;
assign w1126 = 0;
assign w1127 = x5 ? w1153 : w1152;
assign w1128 = 1;
assign w1129 = x14 ? w1155 : w1154;
assign w1130 = x1 ? w1157 : w1156;
assign w1131 = x14 ? w1159 : w1158;
assign w1132 = 0;
assign w1133 = x8 ? w1161 : w1160;
assign w1134 = x10 ? w1163 : w1162;
assign w1135 = x5 ? w1165 : w1164;
assign w1136 = 0;
assign w1137 = x5 ? w1167 : w1166;
assign w1138 = x5 ? w1169 : w1168;
assign w1139 = 0;
assign w1140 = 0;
assign w1141 = x4 ? w1171 : w1170;
assign w1142 = 0;
assign w1143 = x5 ? w1173 : w1172;
assign w1144 = 1;
assign w1145 = x13 ? w1175 : w1174;
assign w1146 = x6 ? w1177 : w1176;
assign w1147 = x13 ? w1179 : w1178;
assign w1148 = 0;
assign w1149 = x3 ? w1181 : w1180;
assign w1150 = 0;
assign w1151 = x5 ? w1183 : w1182;
assign w1152 = 0;
assign w1153 = 1;
assign w1154 = 1;
assign w1155 = 0;
assign w1156 = 1;
assign w1157 = 0;
assign w1158 = 0;
assign w1159 = x1 ? w1185 : w1184;
assign w1160 = 0;
assign w1161 = 1;
assign w1162 = 0;
assign w1163 = 1;
assign w1164 = 1;
assign w1165 = 0;
assign w1166 = 0;
assign w1167 = 1;
assign w1168 = 1;
assign w1169 = 0;
assign w1170 = 0;
assign w1171 = 1;
assign w1172 = 0;
assign w1173 = 1;
assign w1174 = 1;
assign w1175 = 0;
assign w1176 = 1;
assign w1177 = 0;
assign w1178 = 0;
assign w1179 = 1;
assign w1180 = 0;
assign w1181 = 1;
assign w1182 = 1;
assign w1183 = 0;
assign w1184 = 0;
assign w1185 = 1;
assign w101 = x0 ? w103 : w102;
assign w102 = x1 ? w105 : w104;
assign w103 = x13 ? w107 : w106;
assign w104 = x2 ? w109 : w108;
assign w105 = x12 ? w1011 : w1010;
assign w106 = x8 ? w1013 : w1012;
assign w107 = x14 ? w1015 : w1014;
assign w108 = x3 ? w1017 : w1016;
assign w109 = x11 ? w1019 : w1018;
assign w1010 = x8 ? w1021 : w1020;
assign w1011 = x13 ? w1023 : w1022;
assign w1012 = x9 ? w1025 : w1024;
assign w1013 = x6 ? w1027 : w1026;
assign w1014 = x8 ? w1029 : w1028;
assign w1015 = x6 ? w1031 : w1030;
assign w1016 = x4 ? w1033 : w1032;
assign w1017 = x10 ? w1035 : w1034;
assign w1018 = x12 ? w1037 : w1036;
assign w1019 = x12 ? w1039 : w1038;
assign w1020 = x13 ? w1041 : w1040;
assign w1021 = x6 ? w1043 : w1042;
assign w1022 = x14 ? w1045 : w1044;
assign w1023 = x6 ? w1047 : w1046;
assign w1024 = x10 ? w1049 : w1048;
assign w1025 = x5 ? w1051 : w1050;
assign w1026 = x5 ? w1053 : w1052;
assign w1027 = x5 ? w1055 : w1054;
assign w1028 = 1;
assign w1029 = x12 ? w1057 : w1056;
assign w1030 = x1 ? w1059 : w1058;
assign w1031 = 0;
assign w1032 = 0;
assign w1033 = x9 ? w1061 : w1060;
assign w1034 = x11 ? w1063 : w1062;
assign w1035 = x6 ? w1065 : w1064;
assign w1036 = 0;
assign w1037 = x13 ? w1067 : w1066;
assign w1038 = 1;
assign w1039 = x6 ? w1069 : w1068;
assign w1040 = 0;
assign w1041 = x14 ? w1071 : w1070;
assign w1042 = 0;
assign w1043 = 1;
assign w1044 = 1;
assign w1045 = x6 ? w1073 : w1072;
assign w1046 = x2 ? w1075 : w1074;
assign w1047 = 0;
assign w1048 = 0;
assign w1049 = x4 ? w1077 : w1076;
assign w1050 = x4 ? w1079 : w1078;
assign w1051 = 1;
assign w1052 = 0;
assign w1053 = 1;
assign w1054 = x14 ? w1081 : w1080;
assign w1055 = 0;
assign w1056 = 1;
assign w1057 = 0;
assign w1058 = 1;
assign w1059 = x12 ? w1083 : w1082;
assign w1060 = 0;
assign w1061 = 1;
assign w1062 = 0;
assign w1063 = 1;
assign w1064 = 1;
assign w1065 = 0;
assign w1066 = 0;
assign w1067 = 1;
assign w1068 = 1;
assign w1069 = 0;
assign w1070 = 0;
assign w1071 = 1;
assign w1072 = 1;
assign w1073 = 0;
assign w1074 = 1;
assign w1075 = 0;
assign w1076 = 0;
assign w1077 = 1;
assign w1078 = 0;
assign w1079 = 1;
assign w1080 = 0;
assign w1081 = 1;
assign w1082 = 0;
assign w1083 = 1;
assign w91 = x1 ? w93 : w92;
assign w92 = x0 ? w95 : w94;
assign w93 = x13 ? w97 : w96;
assign w94 = x2 ? w99 : w98;
assign w95 = x14 ? w911 : w910;
assign w96 = x9 ? w913 : w912;
assign w97 = x15 ? w915 : w914;
assign w98 = x3 ? w917 : w916;
assign w99 = x12 ? w919 : w918;
assign w910 = x9 ? w921 : w920;
assign w911 = x2 ? w923 : w922;
assign w912 = x8 ? w925 : w924;
assign w913 = x3 ? w927 : w926;
assign w914 = x14 ? w929 : w928;
assign w915 = x7 ? w931 : w930;
assign w916 = x4 ? w933 : w932;
assign w917 = x11 ? w935 : w934;
assign w918 = 0;
assign w919 = x13 ? w937 : w936;
assign w920 = 0;
assign w921 = x5 ? w939 : w938;
assign w922 = 1;
assign w923 = x6 ? w941 : w940;
assign w924 = 0;
assign w925 = x6 ? w943 : w942;
assign w926 = x2 ? w945 : w944;
assign w927 = 1;
assign w928 = x7 ? w947 : w946;
assign w929 = x0 ? w949 : w948;
assign w930 = x9 ? w951 : w950;
assign w931 = 0;
assign w932 = 0;
assign w933 = x10 ? w953 : w952;
assign w934 = 0;
assign w935 = x12 ? w955 : w954;
assign w936 = 1;
assign w937 = x7 ? w957 : w956;
assign w938 = 0;
assign w939 = x7 ? w959 : w958;
assign w940 = 1;
assign w941 = 0;
assign w942 = 0;
assign w943 = x14 ? w961 : w960;
assign w944 = x6 ? w963 : w962;
assign w945 = 0;
assign w946 = x9 ? w965 : w964;
assign w947 = 1;
assign w948 = x2 ? w967 : w966;
assign w949 = x2 ? w969 : w968;
assign w950 = x5 ? w971 : w970;
assign w951 = 1;
assign w952 = 0;
assign w953 = 1;
assign w954 = 1;
assign w955 = 0;
assign w956 = 1;
assign w957 = 0;
assign w958 = 1;
assign w959 = 0;
assign w960 = 1;
assign w961 = 0;
assign w962 = 0;
assign w963 = 1;
assign w964 = 1;
assign w965 = 0;
assign w966 = 1;
assign w967 = 0;
assign w968 = 0;
assign w969 = 1;
assign w970 = 1;
assign w971 = 0;
assign w81 = x0 ? w83 : w82;
assign w82 = x9 ? w85 : w84;
assign w83 = x9 ? w87 : w86;
assign w84 = x7 ? w89 : w88;
assign w85 = x6 ? w811 : w810;
assign w86 = x15 ? w813 : w812;
assign w87 = x6 ? w815 : w814;
assign w88 = x2 ? w817 : w816;
assign w89 = x8 ? w819 : w818;
assign w810 = x11 ? w821 : w820;
assign w811 = x7 ? w823 : w822;
assign w812 = x2 ? w825 : w824;
assign w813 = x7 ? w827 : w826;
assign w814 = x11 ? w829 : w828;
assign w815 = x15 ? w831 : w830;
assign w816 = x1 ? w833 : w832;
assign w817 = x13 ? w835 : w834;
assign w818 = x10 ? w837 : w836;
assign w819 = x10 ? w839 : w838;
assign w820 = x5 ? w841 : w840;
assign w821 = x4 ? w843 : w842;
assign w822 = x15 ? w845 : w844;
assign w823 = x8 ? w847 : w846;
assign w824 = x7 ? w849 : w848;
assign w825 = x13 ? w851 : w850;
assign w826 = x6 ? w853 : w852;
assign w827 = x8 ? w855 : w854;
assign w828 = x15 ? w857 : w856;
assign w829 = x8 ? w859 : w858;
assign w830 = x2 ? w861 : w860;
assign w831 = 0;
assign w832 = 0;
assign w833 = x14 ? w863 : w862;
assign w834 = 0;
assign w835 = x15 ? w865 : w864;
assign w836 = 0;
assign w837 = 1;
assign w838 = 1;
assign w839 = 0;
assign w840 = 0;
assign w841 = x10 ? w867 : w866;
assign w842 = 0;
assign w843 = 1;
assign w844 = x2 ? w869 : w868;
assign w845 = 1;
assign w846 = 0;
assign w847 = 1;
assign w848 = 0;
assign w849 = x8 ? w871 : w870;
assign w850 = 0;
assign w851 = 1;
assign w852 = x11 ? w873 : w872;
assign w853 = 1;
assign w854 = x10 ? w875 : w874;
assign w855 = x10 ? w877 : w876;
assign w856 = 0;
assign w857 = 1;
assign w858 = 1;
assign w859 = 0;
assign w860 = 1;
assign w861 = x13 ? w879 : w878;
assign w862 = 0;
assign w863 = 1;
assign w864 = 1;
assign w865 = 0;
assign w866 = 0;
assign w867 = 1;
assign w868 = 1;
assign w869 = 0;
assign w870 = 0;
assign w871 = 1;
assign w872 = 1;
assign w873 = 0;
assign w874 = 1;
assign w875 = 0;
assign w876 = 0;
assign w877 = 1;
assign w878 = 1;
assign w879 = 0;
assign w71 = x1 ? w73 : w72;
assign w72 = x9 ? w75 : w74;
assign w73 = x9 ? w77 : w76;
assign w74 = x3 ? w79 : w78;
assign w75 = x7 ? w711 : w710;
assign w76 = x15 ? w713 : w712;
assign w77 = x7 ? w715 : w714;
assign w78 = x2 ? w717 : w716;
assign w79 = x13 ? w719 : w718;
assign w710 = x11 ? w721 : w720;
assign w711 = x15 ? w723 : w722;
assign w712 = x3 ? w725 : w724;
assign w713 = x7 ? w727 : w726;
assign w714 = x11 ? w729 : w728;
assign w715 = x15 ? w731 : w730;
assign w716 = x4 ? w733 : w732;
assign w717 = x14 ? w735 : w734;
assign w718 = 0;
assign w719 = x15 ? w737 : w736;
assign w720 = x6 ? w739 : w738;
assign w721 = x5 ? w741 : w740;
assign w722 = x3 ? w743 : w742;
assign w723 = 1;
assign w724 = x14 ? w745 : w744;
assign w725 = x13 ? w747 : w746;
assign w726 = x11 ? w749 : w748;
assign w727 = 1;
assign w728 = x15 ? w751 : w750;
assign w729 = x5 ? w753 : w752;
assign w730 = x3 ? w755 : w754;
assign w731 = 0;
assign w732 = 0;
assign w733 = x12 ? w757 : w756;
assign w734 = 0;
assign w735 = 1;
assign w736 = 1;
assign w737 = x7 ? w759 : w758;
assign w738 = 0;
assign w739 = x10 ? w761 : w760;
assign w740 = 0;
assign w741 = 1;
assign w742 = 1;
assign w743 = x13 ? w763 : w762;
assign w744 = 0;
assign w745 = x2 ? w765 : w764;
assign w746 = 0;
assign w747 = 1;
assign w748 = 1;
assign w749 = x5 ? w767 : w766;
assign w750 = 0;
assign w751 = 1;
assign w752 = 0;
assign w753 = x15 ? w769 : w768;
assign w754 = 1;
assign w755 = x13 ? w771 : w770;
assign w756 = 0;
assign w757 = 1;
assign w758 = 1;
assign w759 = 0;
assign w760 = 0;
assign w761 = 1;
assign w762 = 1;
assign w763 = 0;
assign w764 = 0;
assign w765 = 1;
assign w766 = 1;
assign w767 = 0;
assign w768 = 1;
assign w769 = 0;
assign w770 = 1;
assign w771 = 0;
assign w61 = x2 ? w63 : w62;
assign w62 = x11 ? w65 : w64;
assign w63 = x11 ? w67 : w66;
assign w64 = x7 ? w69 : w68;
assign w65 = x6 ? w611 : w610;
assign w66 = x15 ? w613 : w612;
assign w67 = x6 ? w615 : w614;
assign w68 = x3 ? w617 : w616;
assign w69 = x10 ? w619 : w618;
assign w610 = x12 ? w621 : w620;
assign w611 = x7 ? w623 : w622;
assign w612 = x3 ? w625 : w624;
assign w613 = x7 ? w627 : w626;
assign w614 = x15 ? w629 : w628;
assign w615 = x15 ? w631 : w630;
assign w616 = x4 ? w633 : w632;
assign w617 = x14 ? w635 : w634;
assign w618 = 0;
assign w619 = 1;
assign w620 = 0;
assign w621 = x5 ? w637 : w636;
assign w622 = x15 ? w639 : w638;
assign w623 = x10 ? w641 : w640;
assign w624 = x10 ? w643 : w642;
assign w625 = x14 ? w645 : w644;
assign w626 = x6 ? w647 : w646;
assign w627 = x10 ? w649 : w648;
assign w628 = x3 ? w651 : w650;
assign w629 = x12 ? w653 : w652;
assign w630 = x3 ? w655 : w654;
assign w631 = x7 ? w657 : w656;
assign w632 = 0;
assign w633 = x13 ? w659 : w658;
assign w634 = 0;
assign w635 = x15 ? w661 : w660;
assign w636 = 0;
assign w637 = 1;
assign w638 = x3 ? w663 : w662;
assign w639 = 1;
assign w640 = 0;
assign w641 = 1;
assign w642 = 0;
assign w643 = x7 ? w665 : w664;
assign w644 = 0;
assign w645 = x10 ? w667 : w666;
assign w646 = x12 ? w669 : w668;
assign w647 = 1;
assign w648 = 1;
assign w649 = 0;
assign w650 = x10 ? w671 : w670;
assign w651 = 0;
assign w652 = 1;
assign w653 = x5 ? w673 : w672;
assign w654 = 1;
assign w655 = x10 ? w675 : w674;
assign w656 = 0;
assign w657 = x10 ? w677 : w676;
assign w658 = 0;
assign w659 = 1;
assign w660 = 1;
assign w661 = 0;
assign w662 = 1;
assign w663 = 0;
assign w664 = 0;
assign w665 = 1;
assign w666 = 1;
assign w667 = 0;
assign w668 = 1;
assign w669 = 0;
assign w670 = 0;
assign w671 = 1;
assign w672 = 1;
assign w673 = 0;
assign w674 = 1;
assign w675 = 0;
assign w676 = 1;
assign w677 = 0;
assign w51 = x3 ? w53 : w52;
assign w52 = x11 ? w55 : w54;
assign w53 = x11 ? w57 : w56;
assign w54 = x4 ? w59 : w58;
assign w55 = x7 ? w511 : w510;
assign w56 = x15 ? w513 : w512;
assign w57 = x7 ? w515 : w514;
assign w58 = x5 ? w517 : w516;
assign w59 = x14 ? w519 : w518;
assign w510 = x12 ? w521 : w520;
assign w511 = x15 ? w523 : w522;
assign w512 = x4 ? w525 : w524;
assign w513 = x7 ? w527 : w526;
assign w514 = x15 ? w529 : w528;
assign w515 = x15 ? w531 : w530;
assign w516 = x6 ? w533 : w532;
assign w517 = x13 ? w535 : w534;
assign w518 = 0;
assign w519 = x15 ? w537 : w536;
assign w520 = x4 ? w539 : w538;
assign w521 = x6 ? w541 : w540;
assign w522 = x4 ? w543 : w542;
assign w523 = 1;
assign w524 = x5 ? w545 : w544;
assign w525 = x14 ? w547 : w546;
assign w526 = x12 ? w549 : w548;
assign w527 = 1;
assign w528 = x4 ? w551 : w550;
assign w529 = x12 ? w553 : w552;
assign w530 = x4 ? w555 : w554;
assign w531 = 0;
assign w532 = 0;
assign w533 = x12 ? w557 : w556;
assign w534 = 0;
assign w535 = 1;
assign w536 = 1;
assign w537 = x7 ? w559 : w558;
assign w538 = 0;
assign w539 = x14 ? w561 : w560;
assign w540 = x13 ? w563 : w562;
assign w541 = 1;
assign w542 = 1;
assign w543 = x14 ? w565 : w564;
assign w544 = 0;
assign w545 = x13 ? w567 : w566;
assign w546 = x5 ? w569 : w568;
assign w547 = 1;
assign w548 = 1;
assign w549 = x6 ? w571 : w570;
assign w550 = x12 ? w573 : w572;
assign w551 = x14 ? w575 : w574;
assign w552 = 1;
assign w553 = x6 ? w577 : w576;
assign w554 = 1;
assign w555 = x14 ? w579 : w578;
assign w556 = 0;
assign w557 = 1;
assign w558 = 1;
assign w559 = 0;
assign w560 = 0;
assign w561 = 1;
assign w562 = 0;
assign w563 = 1;
assign w564 = 1;
assign w565 = 0;
assign w566 = 0;
assign w567 = 1;
assign w568 = 0;
assign w569 = 1;
assign w570 = 1;
assign w571 = 0;
assign w572 = 0;
assign w573 = 1;
assign w574 = 0;
assign w575 = 1;
assign w576 = 1;
assign w577 = 0;
assign w578 = 1;
assign w579 = 0;
assign w41 = x4 ? w43 : w42;
assign w42 = x12 ? w45 : w44;
assign w43 = x15 ? w47 : w46;
assign w44 = x5 ? w49 : w48;
assign w45 = x7 ? w411 : w410;
assign w46 = x5 ? w413 : w412;
assign w47 = x12 ? w415 : w414;
assign w48 = x6 ? w417 : w416;
assign w49 = x14 ? w419 : w418;
assign w410 = x13 ? w421 : w420;
assign w411 = x5 ? w423 : w422;
assign w412 = x12 ? w425 : w424;
assign w413 = x14 ? w427 : w426;
assign w414 = x13 ? w429 : w428;
assign w415 = x7 ? w431 : w430;
assign w416 = 0;
assign w417 = x13 ? w433 : w432;
assign w418 = x13 ? w435 : w434;
assign w419 = x6 ? w437 : w436;
assign w420 = x5 ? w439 : w438;
assign w421 = x6 ? w441 : w440;
assign w422 = 1;
assign w423 = x14 ? w443 : w442;
assign w424 = x6 ? w445 : w444;
assign w425 = x7 ? w447 : w446;
assign w426 = x6 ? w449 : w448;
assign w427 = x12 ? w451 : w450;
assign w428 = 1;
assign w429 = x6 ? w453 : w452;
assign w430 = x13 ? w455 : w454;
assign w431 = 0;
assign w432 = 0;
assign w433 = 1;
assign w434 = 0;
assign w435 = x6 ? w457 : w456;
assign w436 = 1;
assign w437 = x15 ? w459 : w458;
assign w438 = 0;
assign w439 = x14 ? w461 : w460;
assign w440 = 0;
assign w441 = 1;
assign w442 = 1;
assign w443 = x15 ? w463 : w462;
assign w444 = 0;
assign w445 = x13 ? w465 : w464;
assign w446 = 0;
assign w447 = 1;
assign w448 = 0;
assign w449 = x13 ? w467 : w466;
assign w450 = 1;
assign w451 = x7 ? w469 : w468;
assign w452 = 1;
assign w453 = x7 ? w471 : w470;
assign w454 = 1;
assign w455 = x6 ? w473 : w472;
assign w456 = 0;
assign w457 = 1;
assign w458 = 1;
assign w459 = 0;
assign w460 = 0;
assign w461 = 1;
assign w462 = 0;
assign w463 = 1;
assign w464 = 0;
assign w465 = 1;
assign w466 = 0;
assign w467 = 1;
assign w468 = 1;
assign w469 = 0;
assign w470 = 0;
assign w471 = 1;
assign w472 = 1;
assign w473 = 0;
assign w31 = x5 ? w33 : w32;
assign w32 = x13 ? w35 : w34;
assign w33 = x15 ? w37 : w36;
assign w34 = x6 ? w39 : w38;
assign w35 = x7 ? w311 : w310;
assign w36 = x6 ? w313 : w312;
assign w37 = x13 ? w315 : w314;
assign w38 = 0;
assign w39 = x14 ? w317 : w316;
assign w310 = x6 ? w319 : w318;
assign w311 = x6 ? w321 : w320;
assign w312 = x7 ? w323 : w322;
assign w313 = x14 ? w325 : w324;
assign w314 = x6 ? w327 : w326;
assign w315 = x7 ? w329 : w328;
assign w316 = 0;
assign w317 = x7 ? w331 : w330;
assign w318 = 0;
assign w319 = x14 ? w333 : w332;
assign w320 = 1;
assign w321 = x14 ? w335 : w334;
assign w322 = 0;
assign w323 = x13 ? w337 : w336;
assign w324 = x7 ? w339 : w338;
assign w325 = x7 ? w341 : w340;
assign w326 = 1;
assign w327 = x7 ? w343 : w342;
assign w328 = x6 ? w345 : w344;
assign w329 = 0;
assign w330 = 1;
assign w331 = x15 ? w347 : w346;
assign w332 = 0;
assign w333 = 1;
assign w334 = 1;
assign w335 = x15 ? w349 : w348;
assign w336 = 0;
assign w337 = 1;
assign w338 = 0;
assign w339 = x13 ? w351 : w350;
assign w340 = 1;
assign w341 = x13 ? w353 : w352;
assign w342 = x14 ? w355 : w354;
assign w343 = 1;
assign w344 = 1;
assign w345 = x14 ? w357 : w356;
assign w346 = 1;
assign w347 = 0;
assign w348 = 0;
assign w349 = 1;
assign w350 = 0;
assign w351 = 1;
assign w352 = 1;
assign w353 = 0;
assign w354 = 1;
assign w355 = 0;
assign w356 = 1;
assign w357 = 0;
assign w21 = x6 ? w23 : w22;
assign w22 = x7 ? w25 : w24;
assign w23 = x15 ? w27 : w26;
assign w24 = 0;
assign w25 = x14 ? w29 : w28;
assign w26 = x7 ? w211 : w210;
assign w27 = x7 ? w213 : w212;
assign w28 = 0;
assign w29 = 1;
assign w210 = 0;
assign w211 = x14 ? w215 : w214;
assign w212 = 1;
assign w213 = x14 ? w217 : w216;
assign w214 = 0;
assign w215 = 1;
assign w216 = 1;
assign w217 = 0;
assign w11 = x7 ? w13 : w12;
assign w12 = 0;
assign w13 = x15 ? w15 : w14;
assign w14 = 0;
assign w15 = 1;
assign y16 = w161;
assign y15 = w151;
assign y14 = w141;
assign y13 = w131;
assign y12 = w121;
assign y11 = w111;
assign y10 = w101;
assign y9 = w91;
assign y8 = w81;
assign y7 = w71;
assign y6 = w61;
assign y5 = w51;
assign y4 = w41;
assign y3 = w31;
assign y2 = w21;
assign y1 = w11;
endmodule
